package fifo_pkg;

endpackage : fifo_pkg
