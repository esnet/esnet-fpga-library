module AXI_tb (
    input dummy
);
endmodule
