package xilinx_hbm_pkg;

endpackage : xilinx_hbm_pkg
