package reg_pkg;

    // Specify data value to return where register access fails (e.g. due to decode error)
    parameter int BAD_ACCESS_DATA = 32'hDEADBEEF;

endpackage : reg_pkg
