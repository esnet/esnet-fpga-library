package sar_verif_pkg;

    import sar_reg_verif_pkg::*;
    import db_verif_pkg::*;
    import htable_verif_pkg::*;
    import state_verif_pkg::*;
    import alloc_verif_pkg::*;
    import state_reg_verif_pkg::*;

    `include "sar_reassembly_htable_reg_agent.svh"
    `include "sar_reassembly_cache_reg_agent.svh"
    `include "sar_reassembly_state_check_reg_agent.svh"
    `include "sar_reassembly_state_reg_agent.svh"
    `include "sar_reassembly_reg_agent.svh"

endpackage : sar_verif_pkg
