package mem_verif_pkg;

    import mem_pkg::*;
    
    `include "mem_agent.svh"

endpackage : mem_verif_pkg
