package reg_verif_pkg;

    // Class definitions
    `include "reg_agent.svh"
    `include "reg_blk_agent.svh"

endpackage : reg_verif_pkg
