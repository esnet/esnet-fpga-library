package reg_pkg;

    // Specify data value to return where register access fails (e.g. due to decode error)
    localparam int BAD_ACCESS_DATA = 32'hDEADBEEF;

endpackage : reg_pkg
