// =============================================================================
//  NOTICE: This computer software was prepared by The Regents of the
//  University of California through Lawrence Berkeley National Laboratory
//  and Jonathan Sewter hereinafter the Contractor, under Contract No.
//  DE-AC02-05CH11231 with the Department of Energy (DOE). All rights in the
//  computer software are reserved by DOE on behalf of the United States
//  Government and the Contractor as provided in the Contract. You are
//  authorized to use this computer software for Governmental purposes but it
//  is not to be released or distributed to the public.
//
//  NEITHER THE GOVERNMENT NOR THE CONTRACTOR MAKES ANY WARRANTY, EXPRESS OR
//  IMPLIED, OR ASSUMES ANY LIABILITY FOR THE USE OF THIS SOFTWARE.
//
//  This notice including this sentence must appear on any copies of this
//  computer software.
// =============================================================================
package db_verif_pkg;

    import db_pkg::*;
    import db_reg_verif_pkg::*;
    
    `include "db_req_transaction.svh"
    `include "db_resp_transaction.svh"
    `include "db_driver.svh"
    `include "db_monitor.svh"
    `include "db_model.svh"
    `include "db_scoreboard.svh"
    `include "db_agent.svh"
    `include "db_ctrl_agent.svh"
    `include "db_reg_agent.svh"

endpackage : db_verif_pkg
