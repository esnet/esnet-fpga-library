package axi4s_verif_pkg;

    // Testbench class definitions
    // (declared here to enforce tb_pkg:: namespace for testbench definitions)
    `include "axi4s_transaction.svh"
    `include "axi4s_driver.svh"
    `include "axi4s_monitor.svh"
    `include "axi4s_sample.svh"
    `include "axi4s_component_env.svh"

endpackage : axi4s_verif_pkg
