package axi4l_verif_pkg;

    // Testbench class definitions
    // (declared here to enforce tb_pkg:: namespace for testbench definitions)
    `include "axi4l_reg_agent.svh"

endpackage : axi4l_verif_pkg
