// =============================================================================
//  NOTICE: This computer software was prepared by The Regents of the
//  University of California through Lawrence Berkeley National Laboratory
//  and Jonathan Sewter hereinafter the Contractor, under Contract No.
//  DE-AC02-05CH11231 with the Department of Energy (DOE). All rights in the
//  computer software are reserved by DOE on behalf of the United States
//  Government and the Contractor as provided in the Contract. You are
//  authorized to use this computer software for Governmental purposes but it
//  is not to be released or distributed to the public.
//
//  NEITHER THE GOVERNMENT NOR THE CONTRACTOR MAKES ANY WARRANTY, EXPRESS OR
//  IMPLIED, OR ASSUMES ANY LIABILITY FOR THE USE OF THIS SOFTWARE.
//
//  This notice including this sentence must appear on any copies of this
//  computer software.
// =============================================================================

interface std_event_intf #(
    parameter type MSG_T = logic
) (
    input logic clk
);
    // Signals
    logic  evt;
    MSG_T  msg;

    // Modports
    modport publisher (
        output evt,
        output msg
    );

    modport subscriber (
        input evt,
        input msg
    );

    clocking cb @(posedge clk);
        default input #1step output #1step;
        output evt, msg;
    endclocking

    task idle();
        cb.evt <= 1'b0;
        cb.msg <= '0;
    endtask

    task _wait(input int cycles);
        repeat (cycles) @(cb);
    endtask

    task notify(input MSG_T _msg);
        cb.evt <= 1'b1;
        cb.msg <= _msg;
        @(cb);
        cb.msg <= 1'b0;
        cb.msg <= '0;
    endtask

endinterface : std_event_intf
