package db_verif_pkg;

    import db_pkg::*;
    import db_reg_verif_pkg::*;
    
    `include "db_req_transaction.svh"
    `include "db_resp_transaction.svh"
    `include "db_driver.svh"
    `include "db_monitor.svh"
    `include "db_model.svh"
    `include "db_scoreboard.svh"
    `include "db_agent.svh"
    `include "db_ctrl_agent.svh"
    `include "db_reg_agent.svh"

endpackage : db_verif_pkg
