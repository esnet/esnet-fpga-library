package mem_proxy_verif_pkg;

    import mem_proxy_reg_verif_pkg::*;
    
    `include "mem_proxy_agent.svh"

endpackage : mem_proxy_verif_pkg
