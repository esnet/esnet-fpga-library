localparam GF_ORDER = 16;
localparam SYM_SIZE = $clog2(GF_ORDER);

localparam logic [SYM_SIZE-1:0] GF_LOG_LUT [GF_ORDER] =
    '{ 1,2,4,8,3,6,12,11,5,10,7,14,15,13,9,0 };

localparam logic [SYM_SIZE-1:0] GF_EXP_LUT [GF_ORDER] =
    '{ 15,0,1,4,2,8,5,10,3,14,9,7,6,13,11,12 };

localparam logic [SYM_SIZE-1:0] GF_MUL_LUT [GF_ORDER][GF_ORDER] = '{
    '{ 0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0 },
    '{ 0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15 },
    '{ 0,2,4,6,8,10,12,14,3,1,7,5,11,9,15,13 },
    '{ 0,3,6,5,12,15,10,9,11,8,13,14,7,4,1,2 },
    '{ 0,4,8,12,3,7,11,15,6,2,14,10,5,1,13,9 },
    '{ 0,5,10,15,7,2,13,8,14,11,4,1,9,12,3,6 },
    '{ 0,6,12,10,11,13,7,1,5,3,9,15,14,8,2,4 },
    '{ 0,7,14,9,15,8,1,6,13,10,3,4,2,5,12,11 },
    '{ 0,8,3,11,6,14,5,13,12,4,15,7,10,2,9,1 },
    '{ 0,9,1,8,2,11,3,10,4,13,5,12,6,15,7,14 },
    '{ 0,10,7,13,14,4,9,3,15,5,8,2,1,11,6,12 },
    '{ 0,11,5,14,10,1,15,4,7,12,2,9,13,6,8,3 },
    '{ 0,12,11,7,5,9,14,2,10,6,1,13,15,3,4,8 },
    '{ 0,13,9,4,1,12,8,5,2,15,11,6,3,14,10,7 },
    '{ 0,14,15,1,13,3,2,12,9,7,6,8,4,10,11,5 },
    '{ 0,15,13,2,9,6,4,11,1,14,12,3,8,7,5,10 }
};

localparam logic [SYM_SIZE-1:0] GF_DIV_LUT [GF_ORDER][GF_ORDER] = '{
    '{ 0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0 },
    '{ 0,1,9,14,13,11,7,6,15,2,12,5,10,4,3,8 },
    '{ 0,2,1,15,9,5,14,12,13,4,11,10,7,8,6,3 },
    '{ 0,3,8,1,4,14,9,10,2,6,7,15,13,12,5,11 },
    '{ 0,4,2,13,1,10,15,11,9,8,5,7,14,3,12,6 },
    '{ 0,5,11,3,12,1,8,13,6,10,9,2,4,7,15,14 },
    '{ 0,6,3,2,8,15,1,7,4,12,14,13,9,11,10,5 },
    '{ 0,7,10,12,5,4,6,1,11,14,2,8,3,15,9,13 },
    '{ 0,8,4,9,2,7,13,5,1,3,10,14,15,6,11,12 },
    '{ 0,9,13,7,15,12,10,3,14,1,6,11,5,2,8,4 },
    '{ 0,10,5,6,11,2,3,9,12,7,1,4,8,14,13,15 },
    '{ 0,11,12,8,6,9,4,15,3,5,13,1,2,10,14,7 },
    '{ 0,12,6,4,3,13,2,14,8,11,15,9,1,5,7,10 },
    '{ 0,13,15,10,14,6,5,8,7,9,3,12,11,1,4,2 },
    '{ 0,14,7,11,10,8,12,2,5,15,4,3,6,13,1,9 },
    '{ 0,15,14,5,7,3,11,4,10,13,8,6,12,9,2,1 }
};

localparam logic [SYM_SIZE-1:0] GF_ADD_LUT [GF_ORDER][GF_ORDER] = '{
    '{ 0,1,2,3,4,5,6,7,8,9,10,11,12,13,14,15 },
    '{ 1,0,3,2,5,4,7,6,9,8,11,10,13,12,15,14 },
    '{ 2,3,0,1,6,7,4,5,10,11,8,9,14,15,12,13 },
    '{ 3,2,1,0,7,6,5,4,11,10,9,8,15,14,13,12 },
    '{ 4,5,6,7,0,1,2,3,12,13,14,15,8,9,10,11 },
    '{ 5,4,7,6,1,0,3,2,13,12,15,14,9,8,11,10 },
    '{ 6,7,4,5,2,3,0,1,14,15,12,13,10,11,8,9 },
    '{ 7,6,5,4,3,2,1,0,15,14,13,12,11,10,9,8 },
    '{ 8,9,10,11,12,13,14,15,0,1,2,3,4,5,6,7 },
    '{ 9,8,11,10,13,12,15,14,1,0,3,2,5,4,7,6 },
    '{ 10,11,8,9,14,15,12,13,2,3,0,1,6,7,4,5 },
    '{ 11,10,9,8,15,14,13,12,3,2,1,0,7,6,5,4 },
    '{ 12,13,14,15,8,9,10,11,4,5,6,7,0,1,2,3 },
    '{ 13,12,15,14,9,8,11,10,5,4,7,6,1,0,3,2 },
    '{ 14,15,12,13,10,11,8,9,6,7,4,5,2,3,0,1 },
    '{ 15,14,13,12,11,10,9,8,7,6,5,4,3,2,1,0 }
};

localparam RS_N  = 10;
localparam RS_K  = 8;
localparam RS_2T = 2;

localparam logic [RS_2T:0][SYM_SIZE-1:0] RS_G_POLY = '{ 8,6,1 };

localparam logic [SYM_SIZE-1:0] RS_G_LUT [RS_K][RS_N] = '{
    '{ 1,0,0,0,0,0,0,0,14,5 },
    '{ 0,1,0,0,0,0,0,0,6,9 },
    '{ 0,0,1,0,0,0,0,0,14,4 },
    '{ 0,0,0,1,0,0,0,0,9,13 },
    '{ 0,0,0,0,1,0,0,0,7,8 },
    '{ 0,0,0,0,0,1,0,0,1,1 },
    '{ 0,0,0,0,0,0,1,0,15,5 },
    '{ 0,0,0,0,0,0,0,1,6,8 }
};

localparam NUM_H = 45;

localparam logic [0:NUM_H-1][0:RS_K-1][0:RS_K-1][SYM_SIZE-1:0] RS_H_LUT = '{
    '{
        '{ 15,9,8,8,7,14,6,14 },
        '{ 4,12,12,13,9,5,9,4 },
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 }
    }, '{
        '{ 7,11,10,13,13,6,12,1 },
        '{ 1,0,0,0,0,0,0,0 },
        '{ 13,3,3,14,15,12,15,1 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 }
    }, '{
        '{ 5,8,1,4,12,12,13,9 },
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 10,14,1,11,5,4,5,14 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 }
    }, '{
        '{ 15,6,1,15,9,8,8,7 },
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 10,14,1,11,5,4,5,14 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 }
    }, '{
        '{ 6,4,7,6,4,3,5,5 },
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 4,3,5,5,2,7,2,3 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 }
    }, '{
        '{ 14,2,13,12,2,13,1,3 },
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 2,8,11,11,9,10,1,8 },
        '{ 0,0,0,0,0,1,0,0 }
    }, '{
        '{ 8,9,3,2,10,3,2,8 },
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 },
        '{ 11,10,13,13,6,12,12,10 }
    }, '{
        '{ 12,10,6,7,11,1,7,11 },
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 },
        '{ 0,0,0,0,0,0,1,0 }
    }, '{
        '{ 10,1,8,9,3,2,10,3 },
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 },
        '{ 0,0,0,0,0,0,1,0 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 6,15,9,8,8,7,14,6 },
        '{ 8,4,12,12,13,9,5,9 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 11,7,11,10,13,13,6,12 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 2,13,3,3,14,15,12,15 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 8,5,8,1,4,12,12,13 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 15,10,14,1,11,5,4,5 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 7,15,6,1,15,9,8,8 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 15,10,14,1,11,5,4,5 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 3,6,4,7,6,4,3,5 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 6,4,3,5,5,2,7,2 },
        '{ 0,0,0,0,0,1,0,0 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 15,14,2,13,12,2,13,1 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 },
        '{ 3,2,8,11,11,9,10,1 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 10,8,9,3,2,10,3,2 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 },
        '{ 0,0,0,0,0,0,1,0 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 12,12,10,6,7,11,1,7 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 },
        '{ 0,0,0,0,0,0,1,0 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 15,6,15,9,8,8,7,14 },
        '{ 5,8,4,12,12,13,9,5 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 7,11,7,11,10,13,13,6 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 12,2,13,3,3,14,15,12 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 13,8,5,8,1,4,12,12 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 4,15,10,14,1,11,5,4 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 9,7,15,6,1,15,9,8 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 4,15,10,14,1,11,5,4 },
        '{ 0,0,0,0,0,1,0,0 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 2,3,6,4,7,6,4,3 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 },
        '{ 7,6,4,3,5,5,2,7 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 12,15,14,2,13,12,2,13 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 },
        '{ 0,0,0,0,0,0,1,0 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 1,10,8,9,3,2,10,3 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 },
        '{ 0,0,0,0,0,0,1,0 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 1,15,6,15,9,8,8,7 },
        '{ 1,5,8,4,12,12,13,9 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 6,7,11,7,11,10,13,13 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 13,12,2,13,3,3,14,15 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 4,13,8,5,8,1,4,12 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 10,4,15,10,14,1,11,5 },
        '{ 0,0,0,0,0,1,0,0 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 14,9,7,15,6,1,15,9 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 },
        '{ 10,4,15,10,14,1,11,5 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 7,2,3,6,4,7,6,4 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 },
        '{ 0,0,0,0,0,0,1,0 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 15,12,15,14,2,13,12,2 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 },
        '{ 0,0,0,0,0,0,1,0 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 7,1,15,6,15,9,8,8 },
        '{ 8,1,5,8,4,12,12,13 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 10,6,7,11,7,11,10,13 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 2,13,12,2,13,3,3,14 },
        '{ 0,0,0,0,0,1,0,0 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 9,4,13,8,5,8,1,4 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 },
        '{ 15,10,4,15,10,14,1,11 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 6,14,9,7,15,6,1,15 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 },
        '{ 0,0,0,0,0,0,1,0 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 2,7,2,3,6,4,7,6 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 },
        '{ 0,0,0,0,0,0,1,0 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 9,7,1,15,6,15,9,8 },
        '{ 13,8,1,5,8,4,12,12 },
        '{ 0,0,0,0,0,1,0,0 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 12,10,6,7,11,7,11,10 },
        '{ 0,0,0,0,0,1,0,0 },
        '{ 14,2,13,12,2,13,3,3 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 5,9,4,13,8,5,8,1 },
        '{ 0,0,0,0,0,1,0,0 },
        '{ 0,0,0,0,0,0,1,0 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 14,6,14,9,7,15,6,1 },
        '{ 0,0,0,0,0,1,0,0 },
        '{ 0,0,0,0,0,0,1,0 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 },
        '{ 14,9,7,1,15,6,15,9 },
        '{ 4,13,8,1,5,8,4,12 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 },
        '{ 1,12,10,6,7,11,7,11 },
        '{ 0,0,0,0,0,0,1,0 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 },
        '{ 9,5,9,4,13,8,5,8 },
        '{ 0,0,0,0,0,0,1,0 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 },
        '{ 0,0,0,0,0,0,1,0 },
        '{ 6,14,9,7,1,15,6,15 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 },
        '{ 0,0,0,0,0,0,1,0 },
        '{ 12,1,12,10,6,7,11,7 }
    }, '{
        '{ 1,0,0,0,0,0,0,0 },
        '{ 0,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,0 },
        '{ 0,0,0,0,0,0,1,0 },
        '{ 0,0,0,0,0,0,0,1 }
    }
};

localparam logic [0:NUM_H-1][0:RS_N-1] RS_ERR_LOC_LUT = '{
        '{ 1,1,0,0,0,0,0,0,0,0 },
        '{ 1,0,1,0,0,0,0,0,0,0 },
        '{ 1,0,0,1,0,0,0,0,0,0 },
        '{ 1,0,0,0,1,0,0,0,0,0 },
        '{ 1,0,0,0,0,1,0,0,0,0 },
        '{ 1,0,0,0,0,0,1,0,0,0 },
        '{ 1,0,0,0,0,0,0,1,0,0 },
        '{ 1,0,0,0,0,0,0,0,1,0 },
        '{ 1,0,0,0,0,0,0,0,0,1 },
        '{ 0,1,1,0,0,0,0,0,0,0 },
        '{ 0,1,0,1,0,0,0,0,0,0 },
        '{ 0,1,0,0,1,0,0,0,0,0 },
        '{ 0,1,0,0,0,1,0,0,0,0 },
        '{ 0,1,0,0,0,0,1,0,0,0 },
        '{ 0,1,0,0,0,0,0,1,0,0 },
        '{ 0,1,0,0,0,0,0,0,1,0 },
        '{ 0,1,0,0,0,0,0,0,0,1 },
        '{ 0,0,1,1,0,0,0,0,0,0 },
        '{ 0,0,1,0,1,0,0,0,0,0 },
        '{ 0,0,1,0,0,1,0,0,0,0 },
        '{ 0,0,1,0,0,0,1,0,0,0 },
        '{ 0,0,1,0,0,0,0,1,0,0 },
        '{ 0,0,1,0,0,0,0,0,1,0 },
        '{ 0,0,1,0,0,0,0,0,0,1 },
        '{ 0,0,0,1,1,0,0,0,0,0 },
        '{ 0,0,0,1,0,1,0,0,0,0 },
        '{ 0,0,0,1,0,0,1,0,0,0 },
        '{ 0,0,0,1,0,0,0,1,0,0 },
        '{ 0,0,0,1,0,0,0,0,1,0 },
        '{ 0,0,0,1,0,0,0,0,0,1 },
        '{ 0,0,0,0,1,1,0,0,0,0 },
        '{ 0,0,0,0,1,0,1,0,0,0 },
        '{ 0,0,0,0,1,0,0,1,0,0 },
        '{ 0,0,0,0,1,0,0,0,1,0 },
        '{ 0,0,0,0,1,0,0,0,0,1 },
        '{ 0,0,0,0,0,1,1,0,0,0 },
        '{ 0,0,0,0,0,1,0,1,0,0 },
        '{ 0,0,0,0,0,1,0,0,1,0 },
        '{ 0,0,0,0,0,1,0,0,0,1 },
        '{ 0,0,0,0,0,0,1,1,0,0 },
        '{ 0,0,0,0,0,0,1,0,1,0 },
        '{ 0,0,0,0,0,0,1,0,0,1 },
        '{ 0,0,0,0,0,0,0,1,1,0 },
        '{ 0,0,0,0,0,0,0,1,0,1 },
        '{ 0,0,0,0,0,0,0,0,1,1 }
};
