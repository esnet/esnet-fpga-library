package timer_verif_pkg;

    import timer_reg_verif_pkg::*;

    // Testbench class definitions
    // (declared here to enforce tb_pkg:: namespace for testbench definitions)
    `include "timer_expiry_reg_agent.svh"

endpackage : timer_verif_pkg
