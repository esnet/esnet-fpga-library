package packet_verif_pkg;
    `include "packet.svh"
    `include "packet_raw.svh"
    `include "packet_eth.svh"
    `include "packet_transaction.svh"

endpackage : packet_verif_pkg

