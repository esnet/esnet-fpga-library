`include "svunit_defines.svh"

// (Failsafe) timeout
`define SVUNIT_TIMEOUT 500us

module rs_decode_unit_test;

    import svunit_pkg::svunit_testcase;
    import std_verif_pkg::*;
    import bus_verif_pkg::*;
    import tb_pkg::*;
    import fec_pkg::*;

    string name = $sformatf("rs_decode_ut");

    svunit_testcase svunit_ut;

    //===================================
    // Parameters
    //===================================
    localparam int DATA_IN_WID = RS_K * SYM_SIZE;

    //===================================
    // Derived parameters
    //===================================

    //===================================
    // Typedefs
    //===================================
    typedef logic [RS_K -1:0][SYM_SIZE-1:0] DATA_IN_T;
    typedef logic [RS_2T-1:0][SYM_SIZE-1:0] PARITY_OUT_T;

    //===================================
    // DUTs (rs_encode -> inject_error -> rs_decode_h_select -> rs_decode)
    //===================================
    logic clk;
    logic srst;

    DATA_IN_T  data_in;
    logic      data_in_valid;
    logic      data_in_ready;

    DATA_IN_T  data_out;
    PARITY_OUT_T parity_out;
    logic      data_out_valid;
    logic      data_out_ready;

    rs_encode DUT0 (.*);


    DATA_IN_T  hsel_data_in = '0;
    logic      [$clog2(NUM_H)-1:0] hsel_err_loc = '0;

    always @(negedge clk) if (data_out_valid)
        inject_error (
            .data_in   (data_out),
            .parity_in (parity_out),
            .data_out  (hsel_data_in),
            .err_loc   (hsel_err_loc) );


    DATA_IN_T  hsel_data_out;
    logic      [RS_K-1:0][RS_K-1:0][SYM_SIZE-1:0] hsel_h_matrix;
    logic      [RS_N-1:0] hsel_err_loc_sel;
    logic      hsel_valid;
    logic      hsel_ready;

    rs_decode_h_select DUT1 (
        .clk            (clk),
        .srst           (srst),

        .data_in        (hsel_data_in),
        .err_loc        (hsel_err_loc),
        .data_in_valid  (data_out_valid),
        .data_in_ready  (data_out_ready),

        .data_out       (hsel_data_out),
        .h_matrix       (hsel_h_matrix),
        .err_loc_sel    (hsel_err_loc_sel),
        .data_out_valid (hsel_valid),
        .data_out_ready (hsel_ready)
    );


    DATA_IN_T  rsd_data_out;
    logic      rsd_valid;
    logic      rsd_ready;

    rs_decode DUT2 (
        .clk            (clk),
        .srst           (srst),

        .data_in        (hsel_data_out),
        .h_matrix       (hsel_h_matrix),
        .err_loc_sel    (hsel_err_loc_sel),
        .data_in_valid  (hsel_valid),
        .data_in_ready  (hsel_ready),

        .data_out       (rsd_data_out),
        .data_out_valid (rsd_valid),
        .data_out_ready (rsd_ready)
    );


    function void inject_error (
        input  DATA_IN_T     data_in,
        input  PARITY_OUT_T  parity_in,

        output DATA_IN_T     data_out,
        output [$clog2(NUM_H)-1:0]  err_loc
    );

        logic [RS_N-1:0][SYM_SIZE-1:0] data;
        int num_errors;

        err_loc = $urandom % NUM_H;

        // delete error locations and compress data_out
        data = {parity_in, data_in};
        num_errors=0;
        for (int i=0; i<RS_N; i++)
            if (RS_ERR_LOC_LUT[err_loc][i] == 1'b0) data[i-num_errors] = data[i];
            else num_errors++;

        data_out = data[RS_K-1:0];
        //$display ("err_loc = %d, data_out = %h", err_loc, data_out);

    endfunction // inject_error


    //===================================
    // Testbench
    //===================================
    rs_decode_tb_env #(1, DATA_IN_T) env;  // NUM_THREADS=1

    bus_intf #(DATA_IN_WID) wr_if (.clk);
    bus_intf #(DATA_IN_WID) rd_if (.clk);

    std_reset_intf reset_if (.clk);

    // Assign reset interface
    assign srst = reset_if.reset;

    initial reset_if.ready = 1'b0;
    always @(posedge clk) reset_if.ready <= ~srst;

    // Assign data interfaces
    assign data_in_valid  = wr_if.valid;
    assign data_in        = wr_if.data;
    assign wr_if.ready    = data_in_ready;

    assign rsd_ready      = rd_if.ready;
    assign rd_if.data     = rsd_data_out;
    assign rd_if.valid    = rsd_valid;

    // Assign clock (100MHz)
    `SVUNIT_CLK_GEN(clk, 5ns);

    //===================================
    // Build
    //===================================
    function void build();
        svunit_ut = new(name);

        // Create testbench environment
        env = new("rs_encode_tb_env", reset_if, wr_if, rd_if);
        env.build();
        env.set_debug_level(1);

    endfunction

    //===================================
    // Setup for running the Unit Tests
    //===================================
    task setup();
        svunit_ut.setup();
        env.run();

        #50ns;

    endtask

    //===================================
    // Here we deconstruct anything we
    // need after running the Unit Tests
    //===================================
    task teardown();
        svunit_ut.teardown();

    endtask

    //===================================
    // All tests are defined between the
    // SVUNIT_TESTS_BEGIN/END macros
    //
    // Each individual test must be
    // defined between `SVTEST(_NAME_)
    // `SVTEST_END
    //
    // i.e.
    //   `SVTEST(mytest)
    //     <test code>
    //   `SVTEST_END
    //===================================

    std_verif_pkg::raw_transaction#(DATA_IN_T) transaction_in;

    DATA_IN_T transaction_in_data;
    initial begin
        transaction_in_data[0]=1;
        transaction_in_data[1]=2;
        transaction_in_data[2]=3;
        transaction_in_data[3]=4;
        transaction_in_data[4]=5;
        transaction_in_data[5]=6;
        transaction_in_data[6]=7;
        transaction_in_data[7]=8;
    end

    bit rx_done=0;
    string msg;


    `SVUNIT_TESTS_BEGIN

        `SVTEST(reset)
        `SVTEST_END

        `SVTEST(basic_sanity)
            int N=500;

            for (int i=0; i<N; i++) begin
                // Send transaction
                for (int j=0; j<RS_N; j++) transaction_in_data[j] = $urandom;
                transaction_in = new("transaction_in", transaction_in_data);
                env.inbox.put(transaction_in);
            end

            fork
                #10us if (!rx_done) `INFO("TIMEOUT! waiting for rx packets...");

                while (!rx_done) #100ns if (env.scoreboard.exp_pending()==0) rx_done=1;
            join_any
	      
            #100ns;
            `FAIL_IF_LOG( env.scoreboard.report(msg) > 0, msg );
            `FAIL_UNLESS_EQUAL( env.scoreboard.got_matched(), N );
        `SVTEST_END

    `SVUNIT_TESTS_END

endmodule : rs_decode_unit_test
