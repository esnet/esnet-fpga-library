package tb_pkg;

    `include "rs_encode_tb_env.svh"
    `include "rs_decode_tb_env.svh"

endpackage : tb_pkg
