    function void set_backpressure(input int __backpressure);
        __BACKPRESSURE = __backpressure;
    endfunction
