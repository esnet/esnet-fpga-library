package std_pkg;

endpackage : std_pkg

