package fec_verif_pkg;

    `include "rs_model.svh"

endpackage : fec_verif_pkg
