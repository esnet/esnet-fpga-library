module Packet_tb (
    input dummy
);
endmodule
