package axi4s_verif_pkg;

    // Verif class definitions
    `include "axi4s_transaction.svh"
    `include "axi4s_driver.svh"
    `include "axi4s_monitor.svh"
    `include "axi4s_sample.svh"
    `include "axi4s_component_env.svh"

endpackage : axi4s_verif_pkg
