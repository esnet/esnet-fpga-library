package arb_pkg;

    // -----------------------------
    // Typedefs
    // -----------------------------
    typedef enum {
        RR,
        WCRR
    } arb_rr_mode_t;

endpackage : arb_pkg
