package tb_pkg;
    import std_verif_pkg::*;
    import axi4l_verif_pkg::*;
    import state_verif_pkg::*;

    // Testbench class definitions
    // (declared here to enforce tb_pkg:: namespace for testbench definitions)
    `include "tb_env.svh"

endpackage : tb_pkg
