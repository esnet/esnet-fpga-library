package fifo_pkg;

    // -----------------------------
    // Typedefs
    // -----------------------------
    typedef enum {
        OPT_MODE_TIMING,
        OPT_MODE_LATENCY
    } opt_mode_t;

endpackage : fifo_pkg
