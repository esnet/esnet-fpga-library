// -----------------------------------------------------------------------------
// axi4s_pkt_discard_ovfl is used to discard the full ingress packet when an axi4s 
// data transaction fails due fifo overflow.   This component should be used on 
// any axi4s interface that ignores the tready flow control signal. 
// axi4s_pkt_discard_ovfl is a synchronous component which employs a memory sized to
// buffer up to 3 max packets.
// -----------------------------------------------------------------------------

module axi4s_pkt_discard_ovfl
   import axi4s_pkg::*;
#(
   parameter int MAX_PKT_LEN = 9100, // max number of bytes per packet.
   parameter bit DROP_ERRORED = 0    // when 1, drop 'errored' packets, where error status is carried in lsb of axi4s_in.TUSER
)  (
   axi4s_intf.rx   axi4s_in,
   axi4s_intf.tx   axi4s_out
);

   // axi4s_in interface params
   localparam int DATA_BYTE_WID = axi4s_in.DATA_BYTE_WID;
   localparam int TID_WID       = axi4s_in.TID_WID;
   localparam int TDEST_WID     = axi4s_in.TDEST_WID;
   localparam int TUSER_WID     = axi4s_in.TUSER_WID;

   // Parameter check
   initial begin
       std_pkg::param_check(axi4s_out.DATA_BYTE_WID, DATA_BYTE_WID, "axi4s_out.DATA_BYTE_WID");
       std_pkg::param_check(axi4s_out.TID_WID,       TID_WID,       "axi4s_out.TID_WID");
       std_pkg::param_check(axi4s_out.TDEST_WID,     TDEST_WID,     "axi4s_out.TDEST_WID");
       std_pkg::param_check(axi4s_out.TUSER_WID,     TUSER_WID,     "axi4s_out.TUSER_WID");
   end

   // fifo params
   localparam int MAX_PKT_WRDS = $ceil($itor(MAX_PKT_LEN) / $itor(DATA_BYTE_WID));
   localparam int FIFO_DEPTH   = MAX_PKT_WRDS * 3;  // depth supports 3 max pkts.
   localparam int ADDR_WID     = $clog2(FIFO_DEPTH);

   // error detection signals
   logic [TUSER_WID-1:0] tuser_in;
   logic pkt_error;

   // ovfl discard signals
   logic [ADDR_WID:0] sop_ptr;
   logic              discard;
   logic              tx_pending;

   // fifo context signals
   logic [ADDR_WID:0] wr_ptr, wr_ptr_p, wr_ptr_nxt;
   logic [ADDR_WID:0] rd_ptr;
   logic              rd_req;

   logic [ADDR_WID:0] fill_level;
   logic              almost_full;
   logic              ovfl;
   logic              empty;



   // _axis4s_in signal assignments.
   axi4s_intf #(.DATA_BYTE_WID(DATA_BYTE_WID), .TID_WID(TID_WID), .TDEST_WID(TDEST_WID), .TUSER_WID(TUSER_WID)) 
              _axi4s_in (.aclk(axi4s_in.aclk), .aresetn(axi4s_in.aresetn));

   assign _axi4s_in.tvalid  = axi4s_in.tvalid;
   assign _axi4s_in.tdata   = axi4s_in.tdata;
   assign _axi4s_in.tkeep   = axi4s_in.tkeep;
   assign _axi4s_in.tdest   = axi4s_in.tdest;
   assign _axi4s_in.tid     = axi4s_in.tid;
   assign _axi4s_in.tlast   = axi4s_in.tlast;
   assign _axi4s_in.tuser   = axi4s_in.tuser;

   assign axi4s_in.tready = _axi4s_in.tready && !(discard || ovfl);


   // ---- error detection logic ----
   assign tuser_in = axi4s_in.tuser;
   assign pkt_error = DROP_ERRORED && tuser_in[0];


   // ---- ovfl discard logic ----
   always @(posedge axi4s_in.aclk)
      if (!axi4s_in.aresetn) begin
         sop_ptr <= 0;
         discard <= 0;
      end else begin
         if (axi4s_in.tready && axi4s_in.tvalid && axi4s_in.tlast && !pkt_error) sop_ptr <= wr_ptr_nxt; // save last sop pointer.

         // if discard is asserted, deassert discard at the end of the inbound packet.
	 // else assert discard signal when fifo overflow occurs.
         if (discard && axi4s_in.tvalid && axi4s_in.tlast) discard <= 1'b0;
         else if (ovfl) discard <= 1'b1;
      end


   // ---- write context logic ----
   assign wr_ptr_nxt = wr_ptr + 1;

   always @(posedge axi4s_in.aclk)
      if (!axi4s_in.aresetn) wr_ptr <= '0;   
      else if (axi4s_in.tvalid) begin
	 // restore sop pointer when tlast is asserted and a discard is in progress or a pkt error is detected.
	 // otherwise increment pointer for each valid transfer.
         if (axi4s_in.tlast && (discard || pkt_error))  wr_ptr <= sop_ptr;
         else if (axi4s_in.tready)                      wr_ptr <= wr_ptr_nxt;
      end

   // assert almost_full when there is only FIFO space for one more ingress packet.
   assign fill_level  = wr_ptr-rd_ptr;
   assign almost_full = fill_level > (FIFO_DEPTH-MAX_PKT_WRDS);

   // assert fifo_overflow if almost_full is asserted when new packet arrives i.e. tvalid && sop.
   assign ovfl = almost_full && axi4s_in.tvalid && axi4s_in.sop;





   // ---- pkt buffer instantiation ----
   axi4s_pkt_buffer #(
      .ADDR_WID (ADDR_WID)
   ) axi4s_pkt_buffer_0 (
      .axi4s_in    (_axi4s_in),
      .axi4s_out   (axi4s_out),
      .rd_req      (rd_req),
      .rd_ptr      (rd_ptr),
      .wr_ptr      (wr_ptr),
      .wr_ptr_p    (wr_ptr_p)
   );




   // ---- read context logic ----
   assign rd_req  = axi4s_out.tready && !empty && !tx_pending;

   always @(posedge axi4s_out.aclk)
      if (!axi4s_out.aresetn)  rd_ptr <= 0;
      else if (rd_req)         rd_ptr <= rd_ptr + 1;

   // assert tx_pending if rd_ptr reaches sop_ptr.
   // defers transfer until sop is overwritten on tlast, and the full packet is buffered.
   assign tx_pending = (rd_ptr == sop_ptr);

   // assert empty when pipelined wr_ptr equals rd_ptr.
   assign empty = (rd_ptr == wr_ptr_p);

endmodule
