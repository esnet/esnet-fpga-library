package std_verif_pkg;

    // Base classes
    `include "base.svh"
    `include "transaction.svh"
    `include "component.svh"
    `include "agent.svh"
    `include "driver.svh"
    `include "monitor.svh"
    `include "model.svh"
    `include "predictor.svh"
    `include "scoreboard.svh"
    `include "env.svh"

    // Basic implementation classes
    `include "event_scoreboard.svh"

    `include "raw_transaction.svh"
    `include "raw_model.svh"
    `include "raw_predictor.svh"
    `include "raw_scoreboard.svh"

    `include "basic_env.svh"
    `include "component_env.svh"
    `include "component_ctrl_env.svh"

    `include "wire_model.svh"
    `include "wire_env.svh"

endpackage : std_verif_pkg

