package xilinx_vitisnetp4_example_pkg;
    localparam int TDATA_NUM_BYTES = 1;
    localparam int USER_META_DATA_WIDTH = 1;

    import vitis_net_p4_dpi_pkg::*;
    `include "example_design_pkg.sv"

endpackage : xilinx_vitisnetp4_example_pkg
