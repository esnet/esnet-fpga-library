package xilinx_vitisnetp4_verif_pkg;

   `include "xilinx_vitisnetp4_agent.svh"

endpackage : xilinx_vitisnetp4_verif_pkg

