class axi4s_monitor #(
    parameter int DATA_BYTE_WID = 8,
    parameter type TID_T = bit,
    parameter type TDEST_T = bit,
    parameter type TUSER_T = bit
) extends std_verif_pkg::monitor#(axi4s_transaction#(TID_T, TDEST_T, TUSER_T));

    local static const string __CLASS_NAME = "axi4s_verif_pkg::axi4s_monitor";

    localparam int TID_WID = $bits(TID_T);
    localparam int TDEST_WID = $bits(TDEST_T);
    localparam int TUSER_WID = $bits(TUSER_T);

    //===================================
    // Properties
    //===================================
    local int __tpause = 0;
    local int __MAX_PKT_SIZE = 65536;

    //===================================
    // Interfaces
    //===================================
    virtual axi4s_intf #(
        .DATA_BYTE_WID(DATA_BYTE_WID),
        .TID_WID  (TID_WID),
        .TDEST_WID(TDEST_WID),
        .TUSER_WID(TUSER_WID)
    ) axis_vif;

    //===================================
    // Methods
    //===================================
    // Constructor
    function new(input string name="axi4s_monitor");
        super.new(name);
        // WORKAROUND-INIT-PROPS {
        //     Provide/repeat default assignments for all remaining instance properties here.
        //     Works around an apparent object initialization bug (as of Vivado 2024.2)
        //     where properties are not properly allocated when they are not assigned
        //     in the constructor.
        this.__tpause = 0;
        this.__MAX_PKT_SIZE = 65536;
        this.axis_vif = null;
        // } WORKAROUND-INIT-PROPS
    endfunction

    // Destructor
    // [[ implements std_verif_pkg::base.destroy() ]]
    virtual function automatic void destroy();
        axis_vif = null;
        super.destroy();
    endfunction

    // Configure trace output
    // [[ overrides std_verif_pkg::base.trace_msg() ]]
    function automatic void trace_msg(input string msg);
        _trace_msg(msg, __CLASS_NAME);
    endfunction

    // Set tpause value used by monitor (for stalling receive transactions)
    function automatic void set_tpause(input int tpause);
        this.__tpause = tpause;
    endfunction

    // Set/get receive packet size limit
    // (Used as upper bound on number of bytes received in a given transaction
    //  before the simulation is terminated (with $fatal).
    //  Guards against unbounded memory allocation due to protocol errors
    //  during simulation.)
    function void set_max_pkt_size(input int MAX_PKT_SIZE);
        this.__MAX_PKT_SIZE = MAX_PKT_SIZE;
    endfunction

    function int get_max_pkt_size();
        return this.__MAX_PKT_SIZE;
    endfunction

    // Reset monitor
    // [[ overrides std_verif_pkg::monitor._reset() ]]
    virtual protected function automatic void _reset();
        super._reset();
        this.set_tpause(0);
    endfunction

    // Quiesce AXI-S interface
    // [[ implements std_verif_pkg::component._idle() ]]
    virtual protected task _idle();
        super._idle();
        axis_vif.idle_rx();
    endtask

    // Receive transaction (represented as raw byte array with associated metadata)
    task receive_raw(
            output byte    data[],
            output TID_T   id,
            output TDEST_T dest,
            output TUSER_T user,
            input  int     tpause = 0
        );
        byte __data[$];
        // Signals
        bit [DATA_BYTE_WID-1:0][7:0] tdata;
        bit [DATA_BYTE_WID-1:0] tkeep;
        bit tlast = 1'b0;
        bit [TID_WID-1:0] tid;
        bit [TDEST_WID-1:0] tdest;
        bit [TUSER_WID-1:0] tuser;
        int byte_idx = 0;
        int word_idx = 0;
        int byte_cnt = 0;

        debug_msg("receive_raw: Waiting for data...");

        while (!tlast) begin
            axis_vif.receive(tdata, tkeep, tlast, tid, tdest, tuser, tpause);
            trace_msg($sformatf("receive_raw: Received word %0d.", word_idx));

            while (byte_idx < DATA_BYTE_WID) begin
                if (tkeep[byte_idx]) __data.push_back(tdata[byte_idx]);
                byte_idx++;
            end
            byte_cnt += byte_idx;
            if (byte_cnt > this.get_max_pkt_size()) begin
                error_msg($sformatf("Received packet exceeded MAX_PKT_SIZE limit (%0d)", this.get_max_pkt_size()));
                $fatal(2, "Received packet exceeded MAX_PKT_SIZE limit.");
            end
            byte_idx = 0;
            word_idx++;
        end
        debug_msg($sformatf("receive_raw: Done. Received %0d bytes.", byte_cnt));
        data = __data;
        __data.delete();
        id = tid;
        dest = tdest;
        user = tuser;
    endtask


    // Receive AXI-S transaction from AXI-S bus
    // [[ implements std_verif_pkg::monitor._receive() ]]
    protected task _receive(output axi4s_transaction#(TID_T, TDEST_T, TUSER_T) transaction);
        // Signals
        byte data [];
        TID_T tid;
        TDEST_T tdest;
        TUSER_T tuser;

        debug_msg("Waiting for transaction...");

        // Receive transaction
        receive_raw(data, tid, tdest, tuser, this.__tpause);

        // Build Rx AXI-S transaction
        transaction = axi4s_transaction#(TID_T, TDEST_T, TUSER_T)::create_from_bytes(
            "rx_axi4s_transaction",
            data,
            tid,
            tdest,
            tuser
        );

        debug_msg($sformatf("Received %s (%0d bytes).", transaction.get_name(), transaction.size()));
    endtask

    task flush();
        axis_vif.tready = 1'b1;
    endtask

endclass
