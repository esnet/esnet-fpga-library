package fifo_verif_pkg;

    import fifo_reg_verif_pkg::*;

    // Testbench class definitions
    // (declared here to enforce tb_pkg:: namespace for testbench definitions)
    `include "fifo_reg_agent.svh"

endpackage : fifo_verif_pkg
