package reg_proxy_verif_pkg;

    // Imports
    import reg_verif_pkg::*;

    // Class definitions
    `include "reg_proxy_agent.svh"

endpackage : reg_proxy_verif_pkg
