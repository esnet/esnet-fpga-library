package alloc_verif_pkg;

    import alloc_reg_verif_pkg::*;

    // Testbench class definitions
    // (declared here to enforce tb_pkg:: namespace for testbench definitions)
    `include "alloc_reg_agent.svh"

endpackage : alloc_verif_pkg
